module tb_binary_adder_tree;
	reg	[15:0]	A, B, C, D, E;
	reg	clk;
	wire	[15:0]	out;

	binary_adder_tree uut (
		.A(A),
		.B(B),
		.C(C),
		.D(D),
		.E(E),
		.clk(clk),
		.out(out)
	);
	
	initial begin
		clk = 0;
		forever #5 clk = ~clk;
	end
	
	initial begin
		A = 16'b0000_0000_0000_0001; B = 16'b0000_0000_0000_0010; C = 16'b0000_0000_0000_0100; D = 16'b0000_0000_0000_1000; E = 16'b0000_0000_0001_0000;
		#10;
		
		A = 16'b1111_1111_1111_1111; B = 16'b0000_0000_0000_0000; C = 16'b0000_0000_0000_0000; D = 16'b0000_0000_0000_0000; E = 16'b0000_0000_0000_0001;
		#10;
		
		A = 16'b0000_0000_0000_0000; B = 16'b0000_0000_0000_0000; C = 16'b0000_0000_0000_0000; D = 16'b0000_0000_0000_0000; E = 16'b1111_1111_1111_1111;
		#10;
		
		A = 16'b1111_1111_1111_1111; B = 16'b1111_1111_1111_1111; C = 16'b1111_1111_1111_1111; D = 16'b1111_1111_1111_1111; E = 16'b1111_1111_1111_1111;
		#10;
		
		A = 16'b0000_0000_0000_0000; B = 16'b0000_0000_0000_0000; C = 16'b0000_0000_0000_0000; D = 16'b0000_0000_0000_0000; E = 16'b0000_0000_0000_0000;
		#10;
		
		$stop;
	end
	
	initial begin
		$monitor($time," ns: A=%b, B=%b, C=%b, D=%b, E=%b, out=%b", A, B, C, D, E, out);
	end
endmodule