module uart_module (
  input clk,
  input rst,
  input rx,
  output tx,
  input [7:0] data_in,
  output reg [7:0] data_out
);

endmodule