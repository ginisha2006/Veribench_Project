module fft_module (
  input clk,
  input rst,
  input start,
  input [DATA_WIDTH-1:0] data_in,
  output reg [DATA_WIDTH-1:0] data_out,
  output reg done
);

endmodule