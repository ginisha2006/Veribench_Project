timescale 1ns / 1ps
module fft_module #(parameter DATA_WIDTH=16, FFT_POINTS=1024) (
    input clk,
    input rst,
    input start,
    input [DATA_WIDTH-1:0] data_in,
    output [DATA_WIDTH-1:0] data_out,
    output done
);