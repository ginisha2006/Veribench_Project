module fibonacci_gen_tb;

  reg clk;
  reg rst;
  reg start;
  reg [7:0] n;
  wire [7:0] fib;

  fibonacci_gen #(8) dut (clk, rst, start, n, fib);

  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end

  initial begin
    rst = 1;
    #10 rst = 0;
    n = 8;
    start = 1;
    #100 start = 0;
  end

  initial begin
    $monitor("Time: %t, n: %b, fib: %b", $time, n, fib);
  end

endmodule