timescale 1ns / 100ps

module tb_single_port_ram;

parameter WIDTH = 8;
parameter DEPTH = 64;

reg [WIDTH-1:0] data;
reg [DEPTH-1:0] addr;
reg we;
reg clk;
wire [WIDTH-1:0] q;

single_port_ram #(.WIDTH(WIDTH),.DEPTH(DEPTH)) dut (
	.data(data),
	.addr(addr),
	.we(we),
	.clk(clk),
	.q(q)
);

initial begin
	$monitor($time, "data=%b, addr=%d, we=%b, q=%b", data, addr, we, q);
	data = 0;
	addr = 0;
	we = 0;
	clk = 0;
	forever #10 clk = ~clk;
	#20;
	for (int i = 0; i < DEPTH; i++) begin
		data = i;
		addr = i;
		we = 1;
		#10;
		data = 0;
		addr = i;
		we = 0;
		#10;
	end
	data = 0;
	addr = 0;
	we = 0;
	#100;
	data = 255;
	addr = 63;
	we = 1;
	#10;
	data = 0;
	addr = 63;
	we = 0;
	#10;
	data = 127;
	addr = 31;
	we = 1;
	#10;
	data = 0;
	addr = 31;
	we = 0;
	#10;
	data = 0;
	addr = 15;
	we = 1;
	#10;
	data = 0;
	addr = 15;
	we = 0;
	#10;
	data = 0;
	addr = 7;
	we = 1;
	#10;
	data = 0;
	addr = 7;
	we = 0;
	#10;
	data = 0;
	addr = 3;
	we = 1;
	#10;
	data = 0;
	addr = 3;
	we = 0;
	#10;
	data = 0;
	addr = 1;
	we = 1;
	#10;
	data = 0;
	addr = 1;
	we = 0;
	#10;
	data = 0;
	addr = 0;
	we = 1;
	#10;
	data = 0;
	addr = 0;
	we = 0;
	#10;
	data = 0;
	addr = 2;
	we = 1;
	#10;
	data = 0;
	addr = 2;
	we = 0;
	#10;
	data = 0;
	addr = 6;
	we = 1;
	#10;
	data = 0;
	addr = 6;
	we = 0;
	#10;
	data = 0;
	addr = 4;
	we = 1;
	#10;
	data = 0;
	addr = 4;
	we = 0;
	#10;
	data = 0;
	addr = 5;
	we = 1;
	#10;
	data = 0;
	addr = 5;
	we = 0;
	#10;
	data = 0;
	addr = 12;
	we = 1;
	#10;
	data = 0;
	addr = 12;
	we = 0;
	#10;
	data = 0;
	addr = 13;
	we = 1;
	#10;
	data = 0;
	addr = 13;
	we = 0;
	#10;
	data = 0;
	addr = 14;
	we = 1;
	#10;
	data = 0;
	addr = 14;
	we = 0;
	#10;
	data = 0;
	addr = 16;
	we = 1;
	#10;
	data = 0;
	addr = 16;
	we = 0;
	#10;
	data = 0;
	addr = 17;
	we = 1;
	#10;
	data = 0;
	addr = 17;
	we = 0;
	#10;
	data = 0;
	addr = 18;
	we = 1;
	#10;
	data = 0;
	addr = 18;
	we = 0;
	#10;
	data = 0;
	addr = 19;
	we = 1;
	#10;
	data = 0;
	addr = 19;
	we = 0;
	#10;
	data = 0;
	addr = 20;
	we = 1;
	#10;
	data = 0;
	addr = 20;
	we = 0;
	#10;
	data = 0