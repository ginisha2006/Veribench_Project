module single_port_ram (
    input [7:0] data,
    input [5:0] addr,
    input we,
    input clk,
    output reg [7:0] q
);

reg [15:0] ram [31:0];

always @(posedge clk) begin
if (we) ram[addr] <= data;
q <= ram[addr];
end

endmodule