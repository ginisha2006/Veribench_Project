module counter_tb;

  reg clk;
  reg reset;
  reg ena;
  wire [7:0] result;

  counter dut (clk, reset, result, ena);

  initial begin
    clk = 0;
    forever #5 clk = ~clk;
  end

  initial begin
    reset = 1;
    #10 reset = 0;
    #10 ena = 1;
    #100 ena = 0;
  end

  initial begin
    $monitor("Time: %t clk=%b reset=%b ena=%b result=%h", $time, clk, reset, ena, result);
  end

endmodule