module tb_ternary_adder_tree;
    parameter WIDTH = 16;

    reg [WIDTH-1:0] A, B, C, D, E;
    reg CLK;
    wire [WIDTH-1:0] OUT;

    initial begin
        // Initialize inputs
        A = 0; B = 0; C = 0; D = 0; E = 0;
        CLK = 0;
        
        #10 A = 5'd3; B = 5'd4; C = 5'd5; D = 5'd6; E = 5'd7;
        #10 A = 5'd8; B = 5'd9; C = 5'd10; D = 5'd11; E = 5'd12;
        #10 A = 5'd15; B = 5'd16; C = 5'd17; D = 5'd18; E = 5'd19;
        #10 A = 5'd20; B = 5'd21; C = 5'd22; D = 5'd23; E = 5'd24;
        #10 A = 5'd30; B = 5'd31; C = 5'd32; D = 5'd33; E = 5'd34;
        #10 A = 5'd40; B = 5'd41; C = 5'd42; D = 5'd43; E = 5'd44;
        #10 A = 5'd50; B = 5'd51; C = 5'd52; D = 5'd53; E = 5'd54;
        #10 A = 5'd60; B = 5'd61; C = 5'd62; D = 5'd63; E = 5'd64;
        #10 A = 5'd70; B = 5'd71; C = 5'd72; D = 5'd73; E = 5'd74;
        #10 A = 5'd80; B = 5'd81; C = 5'd82; D = 5'd83; E = 5'd84;
        #10 A = 5'd90; B = 5'd91; C = 5'd92; D = 5'd93; E = 5'd94;
        #10 A = 5'd100; B = 5'd101; C = 5'd102; D = 5'd103; E = 5'd104;
        #10 A = 5'd110; B = 5'd111; C = 5'd112; D = 5'd113; E = 5'd114;
        #10 A = 5'd120; B = 5'd121; C = 5'd122; D = 5'd123; E = 5'd124;
        #10 A = 5'd130; B = 5'd131; C = 5'd132; D = 5'd133; E = 5'd134;
        #10 A = 5'd140; B = 5'd141; C = 5'd142; D = 5'd143; E = 5'd144;
        #10 A = 5'd150; B = 5'd151; C = 5'd152; D = 5'd153; E = 5'd154;
        #10 A = 5'd160; B = 5'd161; C = 5'd162; D = 5'd163; E = 5'd164;
        #10 A = 5'd170; B = 5'd171; C = 5'd172; D = 5'd173; E = 5'd174;
        #10 A = 5'd180; B = 5'd181; C = 5'd182; D = 5'd183; E = 5'd184;
        #10 A = 5'd