module tb_binary_adder_tree;
  // Inputs
  reg clk;
  reg [15:0] A, B, C, D, E;
  // Output
  wire [15:0] out;

  // Instantiate the Binary Adder Tree
  binary_adder_tree dut (
    .A(A),
    .B(B),
    .C(C),
    .D(D),
    .E(E),
    .clk(clk),
    .out(out)
  );

  initial begin
    // Clock generation
    clk = 0;
    forever #5 clk = ~clk;
  end

  initial begin
    // Stimulus
    $display("Time	A		B		C		D		E		out");
    #10 A = 16'hAAAA; B = 16'hBBBB; C = 16'hCCCC; D = 16'hDDDD; E = 16'hEEEE; #10;
    A = 16'hFFFF; B = 16'h0000; C = 16'h0000; D = 16'h0000; E = 16'h0000; #10;
    A = 16'h0000; B = 16'h0000; C = 16'h0000; D = 16'h0000; E = 16'hFFFF; #10;
    A = 16'h0000; B = 16'h0000; C = 16'h0000; D = 16'h0000; E = 16'hAAAA; #10;
    $finish;
  end

endmodule