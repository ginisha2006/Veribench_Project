module tb_fibonacci_gen;

  localparam WIDTH = 8;

  reg clk;
  reg rst;
  reg start;
  reg [WIDTH-1:0] n;
  wire [WIDTH-1:0] fib;

  fibonacci_gen #(WIDTH) dut (clk, rst, start, n, fib);

  always #5 clk = ~clk;

  assert (@(posedge clk)
      $past(fib) == (dut.a + dut.b) &&
      $past(dut.a) == dut.b &&
      $past(dut.b) == (dut.a + dut.b));
  assert (@(posedge clk)
      count < n);
  assert (@(posedge clk)
      rst ? (fib == 0) : 1);

endmodule