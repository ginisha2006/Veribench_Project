module tb_digital_filter (
    input clk,
    input rst,
    input [15:0] data_in,
    output reg [15:0] data_out,
    input [15:0] coeff [31:0]
);

wire clk;
reg rst;
reg [15:0] data_in;
wire [15:0] data_out;
reg [15:0] coeff [31:0];

digital_filter #(.DATA_WIDTH(16), .COEFF_WIDTH(16), .NUM_TAPS(32)) dut (
    .clk(clk),
    .rst(rst),
    .data_in(data_in),
    .data_out(data_out),
    .coeff(coeff)
);

always begin
    clk = 1; #5; clk = 0; #5;
end

always @(*) begin assert (@(posedge clk) disable iff (!rst) data_out == 16'b0); end

always @(*) begin assert (@(posedge clk) disable iff (!rst) $stable(data_out)); end

always @(*) begin assert (@(posedge clk) data_in >= 0); end

assert (@(posedge clk) coeff[0] >= 0;
    @(posedge clk) coeff[1] >= 0;
    @(posedge clk) coeff[2] >= 0;
    @(posedge clk) coeff[3] >= 0;
    @(posedge clk) coeff[4] >= 0;
    @(posedge clk) coeff[5] >= 0;
    @(posedge clk) coeff[6] >= 0;
    @(posedge clk) coeff[7] >= 0;
    @(posedge clk) coeff[8] >= 0;
    @(posedge clk) coeff[9] >= 0;
    @(posedge clk) coeff[10] >= 0;
    @(posedge clk) coeff[11] >= 0;
    @(posedge clk) coeff[12] >= 0;
    @(posedge clk) coeff[13] >= 0;
    @(posedge clk) coeff[14] >= 0;
    @(posedge clk) coeff[15] >= 0;
    @(posedge clk) coeff[16] >= 0;
    @(posedge clk) coeff[17] >= 0;
    @(posedge clk) coeff[18] >= 0;
    @(posedge clk) coeff[19] >= 0;
    @(posedge clk) coeff[20] >= 0;
    @(posedge clk) coeff[21] >= 0;
    @(posedge clk) coeff[22] >= 0;
    @(posedge clk) coeff[23] >= 0;
    @(posedge clk) coeff[24] >= 0;
    @(posedge clk) coeff[25] >= 0;
    @(posedge clk) coeff[26] >= 0;
    @(posedge clk) coeff[27] >= 0;
    @(posedge clk) coeff[28] >= 0;
    @(posedge clk) coeff[29] >= 0;
    @(posedge clk) coeff[30] >= 0;
    @(posedge clk) coeff[31] >= 0);

always @(*) begin assert (@(posedge clk) disable iff (!rst) data_out <= 16'd65535); end

always @(*) begin assert (@(posedge clk) disable iff (!rst) data_out >= 16'd0); end

endmodule