module tb_alu_4bit();

  // Inputs
  reg [3:0] a, b;
  reg [2:0] ALU_Sel;
  reg clk;

  // Outputs
  wire [3:0] ALU_Result;
  wire Zero;
  wire Carry;
  wire Overflow;

  // Instantiate the DUT
  alu_4bit UUT (
    .a(a),
    .b(b),
    .ALU_Sel(ALU_Sel),
    .ALU_Result(ALU_Result),
    .Zero(Zero),
    .Carry(Carry),
    .Overflow(Overflow)
  );

  // Clock generation for properties
  initial clk = 0;
  always #5 clk = ~clk;

  // Property: Correct result for addition
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b000) |-> ({Carry, ALU_Result} === a + b)); end end

  // Property: Correct result for subtraction
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b001) |-> ({Carry, ALU_Result} === a - b)); end end

  // Property: Correct result for AND operation
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b010) |-> (ALU_Result === a & b)); end end

  // Property: Correct result for OR operation
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b011) |-> (ALU_Result === a | b)); end end

  // Property: Correct result for XOR operation
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b100) |-> (ALU_Result === a ^ b)); end end

  // Property: Correct result for NOT operation
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b101) |-> (ALU_Result === ~a)); end end

  // Property: Correct result for shift left operation
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b110) |-> (ALU_Result === a << 1)); end end

  // Property: Correct result for shift right operation
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b111) |-> (ALU_Result === a >> 1)); end end

  // Property: Correct zero detection
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Result == 4'b0000) |-> Zero); end end

  // Property: Correct carry detection during addition
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b000) && (a + b >= 16'd16) |-> Carry); end end

  // Property: Correct overflow detection during addition
  always @(*) begin always @(*) begin assert (@(posedge clk) (ALU_Sel == 3'b000) && (a[3] == b[3]) && (ALU_Result[3] != a[3]) |-> Overflow); end end

endmodule