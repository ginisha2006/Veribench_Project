module mod_demod_tb();
    parameter DATA_WIDTH = 16;
    reg clk;
    reg rst;
    reg [DATA_WIDTH-1:0] data_in;
    wire [DATA_WIDTH-1:0] modulated_signal;
    wire [DATA_WIDTH-1:0] demodulated_data;

    initial begin
        $monitor($time, "clk: %b, rst: %b, data_in: %h%b, modulated_signal: %h%b, demodulated_data: %h%b",
            clk, rst, data_in, modulated_signal, demodulated_data);

        clk = 0; rst = 1; data_in = 0;
        #10 rst = 0;
        #20 clk = ~clk;
        repeat (100) begin
            #5 clk = ~clk;
        end

        data_in = 8'hA2;
        #10 data_in = 8'h12;
        #10 data_in = 8'h34;
        #10 data_in = 8'h56;
        #10 data_in = 8'h78;
        #10 data_in = 8'h9a;
        #10 data_in = 8'ha2;
        #10 data_in = 8'hbc;
        #10 data_in = 8'hd4;
        #10 data_in = 8'he6;
        #10 data_in = 8'hf8;
        #10 data_in = 8'hfa;
        #10 data_in = 8'hfc;
        #10 data_in = 8'hd0;
        #10 data_in = 8'he2;
        #10 data_in = 8'h04;
        #10 data_in = 8'h06;
        #10 data_in = 8'h08;
        #10 data_in = 8'h0a;
        #10 data_in = 8'h0c;
        #10 data_in = 8'h0e;
        #10 data_in = 8'h10;
        #10 data_in = 8'h12;
        #10 data_in = 8'h14;
        #10 data_in = 8'h16;
        #10 data_in = 8'h18;
        #10 data_in = 8'h1a;
        #10 data_in = 8'h1c;
        #10 data_in = 8'h1e;
        #10 data_in = 8'h20;
        #10 data_in = 8'h22;
        #10 data_in = 8'h24;
        #10 data_in = 8'h26;
        #10 data_in = 8'h28;
        #10 data_in = 8'h2a;
        #10 data_in = 8'h2c;
        #10 data_in = 8'h2e;
        #10 data_in = 8'h30;
        #10 data_in = 8'h32;
        #10 data_in = 8'h34;
        #10 data_in = 8'h36;
        #10 data_in = 8'h38;
        #10 data_in = 8'h3a;
        #10 data_in = 8'h3c;
        #10 data_in = 8'h3e;
        #10 data_in = 8'h40;
        #10 data_in = 8'h42;
        #10 data_in = 8'h44;
        #10 data_in = 8'h46;
        #10 data_in = 8'h48;
        #10 data_in = 8'h4a;
        #10 data_in = 8'h4c;
        #10 data_in = 8'h4e;
        #10 data_in = 8'h50;
        #10 data_in = 8'h52;
        #10 data_in = 8'h54;
        #10 data_in = 8'h56;
        #10 data_in = 8'h58;
        #10 data_in = 8'h5a;
        #10 data_in = 8'h5c;
        #10 data_in = 8'h5e;
        #10 data_in = 8'h60;
        #10 data_in = 8'h62;
        #10 data_in = 8'h64;
        #10 data_in = 8'h66;
        #10 data_in = 8'h68;
        #10 data_in = 8'h6a;
        #10 data_in = 8'h6c;
        #10 data_in = 8'h6e;
        #10 data_in = 8'h70;
        #10 data_in = 8'h72;
        #10 data_in = 8'h74;
        #10 data_in = 8'h76;
        #10 data_in = 8'h78;