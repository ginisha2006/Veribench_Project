module tb_bcd_to_gray (
    input clk,
    input [3:0] bcd,
    output reg [3:0] gray
);

wire [3:0] dut_gray;

bcd_to_gray #(.BCD_WIDTH(4), .GRAY_WIDTH(4)) dut (
    .bcd(bcd),
    .gray(dut_gray)
);

property p_clk;
    @(posedge clk) disable iff (!reset) (dut_gray == bcd ^ (bcd >> 1));
endproperty

assert property(p_clk);

property p_no_overflow_underflow;
    @(posedge clk) disable iff (!reset) ($countones(bcd) <= 4 && $countones(bcd) >= 0);
endproperty

assert property(p_no_overflow_underflow);

property p_edge_cases;
    @(posedge clk) disable iff (!reset) ((bcd == 4'b0000) |-> (dut_gray == 4'b0000));
    @(posedge clk) disable iff (!reset) ((bcd == 4'b1001) |-> (dut_gray == 4'b1100));
endproperty

assert property(p_edge_cases);

endmodule