module tb_mod_demod;

  parameter DATA_WIDTH = 16;
  reg clk;
  reg rst;
  reg [DATA_WIDTH-1:0] data_in;
  wire [DATA_WIDTH-1:0] modulated_signal;
  wire [DATA_WIDTH-1:0] demodulated_data;

  mod_demod #(
    .DATA_WIDTH(DATA_WIDTH)
  ) dut (
    .clk(clk),
    .rst(rst),
    .data_in(data_in),
    .modulated_signal(modulated_signal),
    .demodulated_data(demodulated_data)
  );

  always #5 clk = ~clk;

  property p_modulation;
    @(posedge clk)
      modulated_signal == data_in ^ {DATA_WIDTH{1'b1}};
  endproperty

  property p_demodulation;
    @(posedge clk)
      demodulated_data == modulated_signal ^ {DATA_WIDTH{1'b1}};
  endproperty

  assert property(p_modulation);
  assert property(p_demodulation);

endmodule