module alu_4bit(
    input [3:0] a,
    input [3:0] b,
    input [2:0] ALU_Sel,
    output reg [3:0] ALU_Result,
    output reg Zero,
    output reg Carry,
    output reg Overflow
);
always @(*) begin
    case(ALU_Sel)
        3'b000: ALU_Result = a & b; // AND
        3'b001: ALU_Result = a | b; // OR
        3'b010: ALU_Result = a ^ b; // XOR
        3'b011: ALU_Result = a + b; // ADD
        3'b100: ALU_Result = a - b; // SUBTRACT
        default: ALU_Result = 4'b0;
    endcase
    
    if(ALU_Result == 4'b0) 
        Zero = 1;
    else 
        Zero = 0;

    case(ALU_Sel)
        3'b011, 3'b100:
            begin
                Carry = a[3]&b[3];
                Overflow = ((a[3]^b[3])&(~(a[3]^ALU_Result[3])));
            end
        default:
            Carry = 0;
            Overflow = 0;
    endcase
end
endmodule